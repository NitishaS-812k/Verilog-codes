// Code your design here
module AND(output Y, input A,B);
  assign Y = A&B;
endmodule