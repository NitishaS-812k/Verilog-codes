// Code your design here
module OR(output Y, input A,B);
  assign Y = A||B;
endmodule