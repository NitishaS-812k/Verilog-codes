// Code your design here
module XOR(output Y, input A,B);
  assign Y = A^B;
endmodule