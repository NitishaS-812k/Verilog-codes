// Code your design here
module XNOR(output Y, input A,B);
  assign Y = ~(A^B);
endmodule